
library ieee;
use ieee.std_logic_1164.all;

architecture top_arch_generic_adder of top is
begin
end architecture;
