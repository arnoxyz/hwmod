use work.vhdldraw_pkg.all;

entity illusions is
end entity;


architecture arch of illusions is
begin
	ouchi : entity work.ouchi;
	concentric : entity work.concentric;
	--checkerboard : entity work.checkerboard;
	--squarecircle : entity work.squarecircle;
end architecture;
