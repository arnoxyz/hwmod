library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

use work.math_pkg.all;
use work.alu_pkg.all;

entity alu_tb is
end entity;

architecture tb of alu_tb is
begin

	-- Instantiate your ALU here

	stimuli : process
	begin
		-- apply your stimulus here
		wait;
	end process;
end architecture;

