library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.sorting_network_pkg.all;

entity sorting_network_tb is

end entity;

architecture arch of sorting_network_tb is

begin

end architecture;
