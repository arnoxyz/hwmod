library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.sorting_network_pkg.all;
use work.util_pkg.all;

architecture top_arch_sorting_network of top is

begin
	
end architecture;
